`ifndef RISC_V_DEF
`define RISC_V_DEF

`define NUM_INT_REG 32
`define XLEN 32 // We use the term XLEN to refer to the width of an integer register in bits (32 or 64)
`define INSTR_OPCODE_LW 32

`endif  // RISC_V_DEF